interface dff_if (input logic clk, input logic rst);
 // logic clk;
  // logic rst;
  logic din;
  logic dout;
endinterface
